* AD8615 SPICE Macro-model
* Description: Amplifier
* Generic Desc: 2.7/5V, CMOS, OP, Fast, RRIO, 1X
* Developed by: VW ADSJ
* Revision History: 08/10/2012 - Updated to new header style
* 2.0 (02/2010)
* Copyright 2010, 2012 by Analog Devices
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model 
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes: VSY=5V, T=25�C
*
* Not Modeled:
*    
* Parameters modeled include: 
*
* END Notes
*
* Node Assignments
*                       noninverting input
*                       |   inverting input
*                       |   |    positive supply
*                       |   |    |   negative supply
*                       |   |    |   |   output
*                       |   |    |   |   |
*                       |   |    |   |   |
.SUBCKT AD8615          1   2   99  50  45
*
* INPUT STAGE
*
M1   4  7  8  8 PIX L=1E-6 W=3.64E-04
M2   6  2  8  8 PIX L=1E-6 W=3.64E-04
M3  14  7 18 18 NIX L=1E-6 W=1.44E-04
M4  16  2 18 18 NIX L=1E-6 W=1.44E-04
RD1  4 50 1.33E+04
RD2  6 50 1.33E+04
RD3 99 14 1.33E+04
RD4 99 16 1.33E+04
C1   4  6 5.95E-14
C2  14 16 5.95E-14
I1  99  8 3.65E-05
I2  18 50 3.65E-05
V1  99  9 -1.087E+01
V2  19 50 1.280E-01
D1   8  9 DX
D2  19 18 DX
EOS  7  1 POLY(4) (73,98) (22,98) (81,98) (83,98) 2.30E-05 1 1 1 1
IOS  1  2 5.00E-14
*
*CMRR
*
E1  72 98 POLY(2) (1,98) (2,98) 0 1.507E-03 1.507E-03
R10 72 73 1.061E+01
R20 73 98 8.842E-02
C10 72 73 1.00E-06
*
* PSRR
*
EPSY 21 98 POLY(1) (99,50) -0.3750E+00 0.750E-01
RPS1 21 22 7.9577E+00
RPS2 22 98 1.061E-02
CPS1 21 22 1.00E-06
*
* VOLTAGE NOISE 
*
VN1 80 98 0
RN1 80 98 16.45E-3
HN  81 98 VN1 4.3E+00
RN2 81 98 1
*
* FLICKER NOISE 
*
DFN 82 98 DNOISE
VFN 82 98 DC 0.6551
HFN 83 98 POLY(1) VFN 1.00E-03 1.00E+00
RFN 83 98 1
*
* INTERNAL VOLTAGE REFERENCE
*
EREF 98  0 POLY(2) (99,0) (50,0) 0 0.5 0.5
GSY  99 50 POLY(1) (99,50) 8.786E-04 1.33E-05
EVP  97 98 (99,50) 0.5
EVN  51 98 (50,99) 0.5
*
* GAIN STAGE
*
G1 98 30 POLY(2) (4,6) (14,16) 0 3.710E-03 3.710E-03
R1 30 98 1.00E+06
RZ 45 31 5.321E+01
CF 30 31 2.975E-10 
V3 32 30 1.50E+00
V4 30 33 1.08E+00
D3 32 97 DX
D4 51 33 DX
*
* OUTPUT STAGE
*
M5  45 46 99 99 POX L=1E-6 W=1.48E-03
M6  45 47 50 50 NOX L=1E-6 W=9.26E-03
EG1 99 46 POLY(1) (98,30) 8.250E-01 1
EG2 47 50 POLY(1) (30,98) 7.000E-01 1

*
* MODELS
*
.MODEL POX PMOS (LEVEL=2,KP=4.00E-05,VTO=-0.7,LAMBDA=0.047,RD=0)
.MODEL NOX NMOS (LEVEL=2,KP=1.00E-05,VTO=+0.6,LAMBDA=0.022,RD=0)
.MODEL PIX PMOS (LEVEL=2,KP=1.50E-05,VTO=-0.5,LAMBDA=0.047)
.MODEL NIX NMOS (LEVEL=2,KP=4.00E-05,VTO=0.5,LAMBDA=0.022)
.MODEL DX D(IS=1E-14,RS=0.1)
.MODEL DNOISE D(IS=1E-14,RS=0,KF=4.83E-11)
*.MODEL DNOISE D(IS=1E-14,RS=0,KF=3.43E-11)
*
*
.ENDS





